----------------------------------------------------------------------------------
-- Company: USAFA
-- Engineer: C3C John Paul Terragnoli
-- 
-- Create Date:    22:56:08 01/22/2014 
-- Design Name: 2's Compliment
-- Module Name:    Lab1_Terragnoli - Behavioral 
-- Project Name: Lab1 
-- Target Devices: 
-- Tool versions: 
-- Description: when given a three bit number in 2's compliment form, it gives the 
-- 2's compliment negation of that three bit number. 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Lab1_Terragnoli is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           C : in  STD_LOGIC;
           X : out  STD_LOGIC;
           Y : out  STD_LOGIC;
           Z : out  STD_LOGIC);
end Lab1_Terragnoli;

architecture Behavioral of Lab1_Terragnoli is
--signal declarations: 
signal D: std_logic;
signal E: std_logic;
signal F: std_logic;
signal H: std_logic;
signal I: std_logic;
signal J: std_logic;
signal K: std_logic;
signal L: std_logic;
signal M: std_logic;
signal N: std_logic;
signal O: std_logic;

begin


end Behavioral;

